module ps(

);

endmodule